module keyexpansion_tb;
reg [0:127] k1;
wire[1407:0] out1;
reg [1407:0] expected_output;  // 기대 출력값

key_expansion ks (k1, out1);


initial begin
$monitor("k= %h , out= %h",k1,out1);
k1=128'h5468617473206D79204B756E67204675;
expected_output = 1408'h5468617473206D79204B756E67204675E232FCF191129188B159E4E6D679A29356082007C71AB18F76435569A03AF7FAD2600DE7157ABC686339E901C3031EFBA11202C9B468BEA1D75157A01452495BB1293B3305418592D210D232C6429B69BD3DC287B87C47156A6C9527AC2E0E4ECC96ED1674EAAA031E863F24B2A8316A8E51EF21FABB4522E43D7A0656954B6CBFE2BF904559FAB2A16480B4F7F1CBD828FDDEF86DA4244ACCC0A4FE3B316F26;
    #10;
    if (out1 === expected_output)
        $display("✅ keyexpansion PASS");
        else
        $display("❌ keyexpansion FAIL");

    $finish;

end
endmodule